tinkerAccess-Hat
R9 5 0 1M
R8 1 7 1k
D4 8 10 DI_1N4001
R2 2 13 150
D5 7 5 DI_1N4001
C1 0 5 1µF IC=0
D1 9 6 DI_1N4001
D2 10 6 DI_1N4001
D3 8 9 DI_1N4001
R4 9 10 1k
R7 1 8 1k
R6 6 0 1k
R1 3 4 330
R3 11 12 300
R5 8 0 1k

*SRC=1N4001;DI_1N4001;Diodes;Si;  50.0V  1.00A  3.00us   Diodes, Inc. diode
.MODEL DI_1N4001 D  ( IS=76.9p RS=42.0m BV=50.0 IBV=5.00u CJO=39.8p  M=0.333 N=1.45 TT=4.32u )

.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END
